`timescale 1 ns / 1 ps

module top (
    input clk,

    output B0_C0,
    output B0_D0,
    output B0_C1,
    output B0_D1,
    output B0_C2,
    output B0_D2,
    output B0_C3,
    output B0_D3,
    output B0_C4,
    output B0_D4,
    output B0_C5,
    output B0_D5,
    output B0_C6,
    output B0_D6,
    output B0_C7,
    output B0_D7,

    output B1_C0,
    output B1_D0,
    output B1_C1,
    output B1_D1,
    output B1_C2,
    output B1_D2,
    output B1_C3,
    output B1_D3,
    output B1_C4,
    output B1_D4,
    output B1_C5,
    output B1_D5,

    output B2_C0,
    output B2_D0,
    output B2_C1,
    output B2_D1,
    output B2_C2,
    output B2_D2,
    output B2_C3,
    output B2_D3,
    output B2_C4,
    output B2_D4,
    output B2_C5,
    output B2_D5,
    output B2_C6,
    output B2_D6,
    output B2_C7,
    output B2_D7,

    output B3_C0,
    output B3_D0,
    output B3_C1,
    output B3_D1,
    output B3_C2,
    output B3_D2,
    output B3_C3,
    output B3_D3,
    output B3_C4,
    output B3_D4,
    output B3_C5,
    output B3_D5
);
    assign B0_C0 = clk;
    assign B0_D0 = clk;
    assign B0_C1 = clk;
    assign B0_D1 = clk;
    assign B0_C2 = clk;
    assign B0_D2 = clk;
    assign B0_C3 = clk;
    assign B0_D3 = clk;
    assign B0_C4 = clk;
    assign B0_D4 = clk;
    assign B0_C5 = clk;
    assign B0_D5 = clk;
    assign B0_C6 = clk;
    assign B0_D6 = clk;
    assign B0_C7 = clk;
    assign B0_D7 = clk;

    assign B1_C0 = clk;
    assign B1_D0 = clk;
    assign B1_C1 = clk;
    assign B1_D1 = clk;
    assign B1_C2 = clk;
    assign B1_D2 = clk;
    assign B1_C3 = clk;
    assign B1_D3 = clk;
    assign B1_C4 = clk;
    assign B1_D4 = clk;
    assign B1_C5 = clk;
    assign B1_D5 = clk;

    assign B2_C0 = clk;
    assign B2_D0 = clk;
    assign B2_C1 = clk;
    assign B2_D1 = clk;
    assign B2_C2 = clk;
    assign B2_D2 = clk;
    assign B2_C3 = clk;
    assign B2_D3 = clk;
    assign B2_C4 = clk;
    assign B2_D4 = clk;
    assign B2_C5 = clk;
    assign B2_D5 = clk;
    assign B2_C6 = clk;
    assign B2_D6 = clk;
    assign B2_C7 = clk;
    assign B2_D7 = clk;

    assign B3_C0 = clk;
    assign B3_D0 = clk;
    assign B3_C1 = clk;
    assign B3_D1 = clk;
    assign B3_C2 = clk;
    assign B3_D2 = clk;
    assign B3_C3 = clk;
    assign B3_D3 = clk;
    assign B3_C4 = clk;
    assign B3_D4 = clk;
    assign B3_C5 = clk;
    assign B3_D5 = clk;
endmodule
